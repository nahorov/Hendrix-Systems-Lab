* ======================================================================
* Fuzz Face — Germanium PNP, positive ground
* Differences from SI version:
*   - Chassis ground (0) is the positive battery terminal.
*   - VNEG sits at −9 V relative to ground.
*   - PNP emitters go to the more positive node (ground).
*
* Matches your Makefile:
*   AC wrdata: frequency, v(in), i(vsig)
*   TRAN wrdata: time, v(out), v(b1), v(c2)
* ======================================================================

************* SUPPLY: DEFINE NEGATIVE RAIL *****************************
Vbat 0 VNEG 9          ; makes VNEG = −9 V (0 is +9 V chassis ground)

************* SOURCE / PICKUP ******************************************
.param VINrms = 0.15
.param VIN    = { VINrms*sqrt(2) }
VSIG IN 0 SIN(0 {VIN} 440) AC 1
Rsrc IN IN1 6k
Cin  IN1 B1 10u

************* PNP CORE *************************************************
* Q1 (PNP): collector pulled toward VNEG via Rc, emitter at ground (0)
Q1 C1 B1 0 QPNP
Rc1 VNEG C1 33k
Re1 0  E1 100

* Bias divider (to put B1 between 0 and VNEG appropriately)
Rb1 0   B1 470k        ; from +9 V (ground) to base
Rb2 B1 VNEG 470k       ; from base to −9 V

* Interstage
Ccou C1 B2 100n
Rbleed B2 0 470k

* Q2 (PNP): output at collector C2
Q2 C2 B2 0 QPNP
Rc2 VNEG C2 8.2k
Re2 0  E2 100
Csh C2 0 100p

* Output (remember ground is the positive rail)
Cout C2 OUT 10u
Rload OUT 0 100k

************* TRANSISTOR MODEL (approx Ge PNP) ************************
.model QPNP PNP (IS=5e-9 BF=120 VAF=60 CJE=20p CJC=12p
+               TF=400p TR=400p RB=200 RE=1 RC=50)

************* ANALYSES *************************************************
.op

* AC: drive is AC 1 at VSIG → measure v(in) and i(vsig)
.ac dec 200 20 20k
.save v(in) i(vsig) v(out)

* TRAN: waveshaping
.tran 0.1ms 200ms 0 1us
.save v(out) v(b1) v(c2) v(in)

* Optional: temperature exploration (your Makefile had a temp driver)
* Uncomment to sweep:
* .step temp 0 50 10

.four 440 v(out)

.end

